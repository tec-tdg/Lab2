module testbenchFullAdder();

logic 
